`ifndef PAC
`define PAC

class Packet;
	rand reg [15:0] PWDATA_i;
endclass

`endif 